INCLUDE ./module_a.spi

.subckt top A B C D
.end
