INCLUDE ./module_b.spi

.subckt AN3 a1 a2 a3
.end
