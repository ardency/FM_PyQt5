.subckt AN3 a3 a2 a1
.end
